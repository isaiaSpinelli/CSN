-------------------------------------------------------------------------------
-- HEIG-VD, Haute Ecole d'Ingenierie et de Gestion du canton de Vaud
-- Institut REDS, Reconfigurable & Embedded Digital Systems
--
-- Fichier      : horloge_top.vhd
--
-- Description  : Comparateur pour les ton et le compteur PWM
--
-- Auteur       : Isaia Spinelli et Gaetan Bacso
-- Date         : 16.01.2020
-- Version      : 1.0

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity horloge_top is
   port(

       );
end horloge_top;

architecture flot_don of horloge_top is

  --internally signals

begin


end horloge_top;
