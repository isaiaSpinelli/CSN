-------------------------------------------------------------------------------
-- HEIG-VD, Haute Ecole d'Ingenierie et de Gestion du canton de Vaud
-- Institut REDS, Reconfigurable & Embedded Digital Systems
--
-- Fichier      : emet_serie_uc.vhd
--
-- Description  : Comparateur pour les ton et le compteur PWM
--
-- Auteur       : Isaia Spinelli et Gaetan Bacso
-- Date         : 16.01.2020
-- Version      : 1.0

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity emet_serie_uc is
   port(

       );
end emet_serie_uc;

architecture flot_don of emet_serie_uc is

  --internally signals

begin


end emet_serie_uc;
